`timescale 1ns / 1ps

module uart_tb_parity_error;
    uart_tb_base #(.TESTCASE_ID(2)) tb();
endmodule
