`timescale 1ns / 1ps

module uart_tb_baud_sweep;
    uart_tb_base #(.TESTCASE_ID(6)) tb();
endmodule
