`timescale 1ns / 1ps

module uart_tb_rx_timeout;
    uart_tb_base #(.TESTCASE_ID(5)) tb();
endmodule
