`timescale 1ns / 1ps

module uart_tb_stop_bits;
    uart_tb_base #(.TESTCASE_ID(3)) tb();
endmodule
