`timescale 1ns / 1ps

module uart_tb_reg_access;
    uart_tb_base #(.TESTCASE_ID(0)) tb();
endmodule
