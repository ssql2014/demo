`timescale 1ns / 1ps

module uart_tb_loopback;
    uart_tb_base #(.TESTCASE_ID(1)) tb();
endmodule
