`timescale 1ns / 1ps

module uart_tb_rx_overflow;
    uart_tb_base #(.TESTCASE_ID(4)) tb();
endmodule
